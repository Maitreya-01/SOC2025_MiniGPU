module tb_Full_adder;

  reg a, b, cin;

  wire sum, cout;

  Full_adder uut (
    .a(a),
    .b(b),
    .cin(cin),
    .sum(sum),
    .cout(cout)
  );

  initial begin
    $display("Time | a b cin | sum cout");
    $monitor("%4t | %b %b  %b  |  %b    %b", $time, a, b, cin, sum, cout);

    a = 0; b = 0; cin = 0; #10;
    a = 0; b = 0; cin = 1; #10;
    a = 0; b = 1; cin = 0; #10;
    a = 0; b = 1; cin = 1; #10;
    a = 1; b = 0; cin = 0; #10;
    a = 1; b = 0; cin = 1; #10;
    a = 1; b = 1; cin = 0; #10;
    a = 1; b = 1; cin = 1; #10;

    $stop;
  end

endmodule
